// ----------------------------------------------------------------------------
// Author:   Konstantin Kurenkov
// Email:    krendkrend@gmail.com
// Create date: 19/10/2022
// FileName: kvt_proj_name_define.sv
//
// Description: Define parameter
//
// ----------------------------------------------------------------------------

`ifndef INC_KVT_proj_name_DEFINE
`define INC_KVT_proj_name_DEFINE

	// `ifndef AXI4_ADDR_WIDTH
	// 	`define AXI4_ADDR_WIDTH 64
	// `endif

	// `ifndef AXI4_DATA_WIDTH
	// 	`define AXI4_DATA_WIDTH 64
	// `endif

`endif // INC_KVT_proj_name_DEFINE