// ----------------------------------------------------------------------------
// Author:   Konstantin Kurenkov
// Email:    krendkrend@gmail.com
// Create date: 19/10/2022
// FileName: kvt_proj_name_env_if.sv
//
// Description: Environment Interface
//
// ----------------------------------------------------------------------------

`ifndef INC_KVT_PROJ_NAME_ENV_IF
`define INC_KVT_PROJ_NAME_ENV_IF

interface kvt_proj_name_env_if();

    //  Clock and the reset.
    // -------------------- //

    // Other Interface
    // -------------------- //

endinterface


`endif // INC_KVT_PROJ_NAME_ENV_IF