// ----------------------------------------------------------------------------
// Author:   Konstantin Kurenkov
// Email:    krendkrend@gmail.com
// FileName: kvt_proj_name_wrapper.sv
// Create date: 18/10/2022
//
// Description: Wrapper for proj_name module
//
// ----------------------------------------------------------------------------

`ifndef INC_KVT_PROJ_NAME_WRAPPER
`define INC_KVT_PROJ_NAME_WRAPPER

module kvt_proj_name_wrapper(kvt_proj_name_env_if proj_name_env_if);

// instance proj_name

endmodule : kvt_proj_name_wrapper

`endif // INC_KVT_PROJ_NAME_WRAPPER