{% extends "_base.sv" %}
{% block body %}

	// `ifndef AXI4_ADDR_WIDTH
	// 	`define AXI4_ADDR_WIDTH 64
	// `endif

	// `ifndef AXI4_DATA_WIDTH
	// 	`define AXI4_DATA_WIDTH 64
	// `endif

{% endblock %}
